// 7-���׸�Ʈ ǥ���� ���� ��� 
// 1�� ���� ��, 0�� ���� ������ ����.
// 8��° ĭ�� ������ ���� ���ϴ� ��(dp)�� �ǹ��ϴµ� ������� ���� ���̹Ƿ� ��� 1�� �Ѵ�.
module seven_segment(input [3:0] digit, output reg [7:0] seg);
    always @(*) begin
        case (digit)
            4'b0000: seg = 8'b11000000; // 0
            4'b0001: seg = 8'b11111001; // 1
            4'b0010: seg = 8'b10100100; // 2
            4'b0011: seg = 8'b10110000; // 3
            4'b0100: seg = 8'b10011001; // 4
            4'b0101: seg = 8'b10010010; // 5
            4'b0110: seg = 8'b10000010; // 6
            4'b0111: seg = 8'b11111000; // 7
            4'b1000: seg = 8'b10000000; // 8
            4'b1001: seg = 8'b10010000; // 9
            default: seg = 8'b11111111; // �̿ܿ� �ٸ� ���ڰ� �Է����� ���� �� ��� off
        endcase
    end
endmodule